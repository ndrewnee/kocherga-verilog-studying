// my_cordic.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module my_cordic (
		input  wire [26:0] a,      //      a.a
		input  wire        areset, // areset.reset
		output wire [9:0]  c,      //      c.c
		input  wire        clk,    //    clk.clk
		output wire [9:0]  s       //      s.s
	);

	my_cordic_CORDIC_0 cordic_0 (
		.clk    (clk),    //    clk.clk
		.areset (areset), // areset.reset
		.a      (a),      //      a.a
		.c      (c),      //      c.c
		.s      (s)       //      s.s
	);

endmodule
